library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


entity ForwardingUnit is
   port(
 
	  -- Outputs:
	  ForwardA 	 : out std_logic_vector(1 downto 0);
	  ForwardB	 : out std_logic_vector(1 downto 0);
	  
	  -- Inputs
	  idexRs 	 : in  std_logic_vector(4 downto 0);
	  idexRt	 : in  std_logic_vector(4 downto 0);
	  
	  exmemRegWrite : in  std_logic;
	  exmemRd	 : in  std_logic_vector(4 downto 0);
	  
	  memwbRegWrite	: in  std_logic;
	  memwbRd	 : in  std_logic_vector(4 downto 0)
   );
end ForwardingUnit;

architecture arqFor of ForwardingUnit is 
	begin

		--ForwardA

			--EX hazard
		ForwardA <= "10" when ((exmemRegWrite = '1' and (exmemRd /= 0))
								and (exmemRd = idexRs)) else	
			--MEM hazard
					"01" when ((memwbRegWrite = '1' and (memwbRd /= 0)) 
								and (memwbRd = idexRs)) else "00";
		
		--ForwardB
		
			--EX hazard
		ForwardB <= "10" when ((exmemRegWrite = '1' and (exmemRd /= 0))
								and (exmemRd = idexRt)) else
				
			--MEM hazard
					"01" when ((memwbRegWrite = '1' and (memwbRd /= 0))
								and (memwbRd = idexRt)) else "00";
		
		

end architecture;